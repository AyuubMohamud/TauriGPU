module gpu_control #(
    parameter WIDTH = 32
)(
    input logic clk_i,

);



endmodule
