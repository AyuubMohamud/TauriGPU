module control_unit #(
    parameter WIDTH = 32
)(
    input wire [7:0] opcode,

);




    
endmodule
