module stencil_buffer #(
    parameter WIDTH = 32;
)(


);


endmodule
