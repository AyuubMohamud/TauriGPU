module decode #(
    parameter WIDTH = 32
)(
    input wire [7:0] opcode,
    output wire [3:0] decoded_output
);


    
endmodule