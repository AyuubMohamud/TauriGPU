module fp_ceil #(
    parameter WIDTH = 24
)(
    input  wire logic [WIDTH - 1:0] a,
    output wire logic [WIDTH - 1:0] result
);

    


endmodule
